----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    20:34:48 12/17/2014 
-- Design Name: 
-- Module Name:    SAVE_subtract - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity SAVE_subtract is
    Port ( input_a : in  STD_LOGIC_VECTOR (31 downto 0);
           input_b : in  STD_LOGIC_VECTOR (31 downto 0);
           output : out  STD_LOGIC_VECTOR (31 downto 0));
end SAVE_subtract;

architecture Behavioral of SAVE_subtract is

begin

LOGIC:
	for i in 0 to 31 generate
	begin
		output(i) <= input_a(i) xor input_b(i);
	end generate;
end Behavioral;

