--------------------------------------------------------------------------------
-- Company: Digilent Inc.
-- Engineer: Mircea Dabacan
--
-- Create Date:    12:04:37 08/18/06
-- Design Name:    Digital Scope
-- Module Name:    BlockRam - Structural
-- Project Name:   
-- Target Device:  
-- Tool versions:  
-- Description:
--   The BlockRam component simply instantiates a 2kX8bit Block RAM,
--   disabling the Set/Reset inputs and Parity bits.
--   The Block Ram content is initialized to all zeros.
--
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
--------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

Library UNISIM;
use UNISIM.vcomponents.all;

entity BlockRam is
	Port ( 
		clkA : in std_logic;
		adrA : in std_logic_vector(10 downto 0);
		busDiA : in std_logic_vector(7 downto 0);
		busDoA : out std_logic_vector(7 downto 0);
		ctlEnA : in std_logic;
		ctlWeA : in std_logic;

		clkB : in std_logic;
		adrB : in std_logic_vector(8 downto 0);
		busDiB : in std_logic_vector(31 downto 0);
		busDoB : out std_logic_vector(31 downto 0);
		ctlEnB : in std_logic;
		ctlWeB : in std_logic);
end BlockRam;

architecture Structural of BlockRam is

	Constant DntCare: std_logic_vector(0 downto 0) := "0";
	Constant DntCare2: std_logic_vector(3 downto 0) := "0000";
	-- DIPA and DIPB are defined as std_logic_vector(0 downto 0)

begin

	-- 512 x 32bit memory block 
	RAMB16_S9_S36_inst : RAMB16_S9_S36
	generic map (
		INIT_A => X"000",  --  Value of output RAM registers on Port A at startup
		INIT_B => X"000",  --  Value of output RAM registers on Port B at startup
		SRVAL_A => X"000", --  Port A output value upon SSR assertion
		SRVAL_B => X"000", --  Port B output value upon SSR assertion
		WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
		WRITE_MODE_B => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
		SIM_COLLISION_CHECK => "ALL",  -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL" 
		INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
		INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
		INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
	port map (
		DOA => busDoA,     -- Port A 8-bit Data Output
		DOB => busDoB,     -- Port B 32-bit Data Output    
		DOPA => open,      -- Port A 1-bit Parity Output
		DOPB => open,      -- Port B 1-bit Parity Output
		ADDRA => adrA,     -- Port A 11-bit Address Input
		ADDRB => adrB,     -- Port B 9-bit Address Input
		CLKA => ClkA,      -- Port A Clock
		CLKB => clkB,      -- Port B Clock
		DIA => busDiA,     -- Port A 8-bit Data Input
		DIB => busDiB,     -- Port B 32-bit Data Input
		DIPA => DntCare,   -- Port A 1-bit parity Input, never used
		DIPB => DntCare2,   -- Port-B 1-bit parity Input, never used
		ENA => ctlEnA,     -- Port A RAM Enable Input
		ENB => ctlEnB,     -- Port B RAM Enable Input
		SSRA => '0',       -- Port A Synchronous Set/Reset Input
		SSRB => '0',       -- Port B Synchronous Set/Reset Input
		WEA => ctlWeA,     -- Port A Write Enable Input
		WEB => ctlWeB      -- Port B Write Enable Input
	);

end Structural;
