----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:16:12 12/05/2014 
-- Design Name: 
-- Module Name:    wdec - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity wdec is
	Port ( size : in  STD_LOGIC_VECTOR (7 downto 0);
		widthv : out  STD_LOGIC_VECTOR (127 downto 0));
end wdec;

architecture Behavioral of wdec is

begin
	with size select
	widthv <= X"00000000000000000000000000000000" when X"00",
		X"80000000000000000000000000000000" when X"01",
		X"C0000000000000000000000000000000" when X"02",
		X"E0000000000000000000000000000000" when X"03",
		X"F0000000000000000000000000000000" when X"04",
		X"F8000000000000000000000000000000" when X"05",
		X"FC000000000000000000000000000000" when X"06",
		X"FE000000000000000000000000000000" when X"07",
		X"FF000000000000000000000000000000" when X"08",
		X"FF800000000000000000000000000000" when X"09",
		X"FFC00000000000000000000000000000" when X"0A",
		X"FFE00000000000000000000000000000" when X"0B",
		X"FFF00000000000000000000000000000" when X"0C",
		X"FFF80000000000000000000000000000" when X"0D",
		X"FFFC0000000000000000000000000000" when X"0E",
		X"FFFE0000000000000000000000000000" when X"0F",
		X"FFFF0000000000000000000000000000" when X"10",
		X"FFFF8000000000000000000000000000" when X"11",
		X"FFFFC000000000000000000000000000" when X"12",
		X"FFFFE000000000000000000000000000" when X"13",
		X"FFFFF000000000000000000000000000" when X"14",
		X"FFFFF800000000000000000000000000" when X"15",
		X"FFFFFC00000000000000000000000000" when X"16",
		X"FFFFFE00000000000000000000000000" when X"17",
		X"FFFFFF00000000000000000000000000" when X"18",
		X"FFFFFF80000000000000000000000000" when X"19",
		X"FFFFFFC0000000000000000000000000" when X"1A",
		X"FFFFFFE0000000000000000000000000" when X"1B",
		X"FFFFFFF0000000000000000000000000" when X"1C",
		X"FFFFFFF8000000000000000000000000" when X"1D",
		X"FFFFFFFC000000000000000000000000" when X"1E",
		X"FFFFFFFE000000000000000000000000" when X"1F",
		X"FFFFFFFF000000000000000000000000" when X"20",
		X"FFFFFFFF800000000000000000000000" when X"21",
		X"FFFFFFFFC00000000000000000000000" when X"22",
		X"FFFFFFFFE00000000000000000000000" when X"23",
		X"FFFFFFFFF00000000000000000000000" when X"24",
		X"FFFFFFFFF80000000000000000000000" when X"25",
		X"FFFFFFFFFC0000000000000000000000" when X"26",
		X"FFFFFFFFFE0000000000000000000000" when X"27",
		X"FFFFFFFFFF0000000000000000000000" when X"28",
		X"FFFFFFFFFF8000000000000000000000" when X"29",
		X"FFFFFFFFFFC000000000000000000000" when X"2A",
		X"FFFFFFFFFFE000000000000000000000" when X"2B",
		X"FFFFFFFFFFF000000000000000000000" when X"2C",
		X"FFFFFFFFFFF800000000000000000000" when X"2D",
		X"FFFFFFFFFFFC00000000000000000000" when X"2E",
		X"FFFFFFFFFFFE00000000000000000000" when X"2F",
		X"FFFFFFFFFFFF00000000000000000000" when X"30",
		X"FFFFFFFFFFFF80000000000000000000" when X"31",
		X"FFFFFFFFFFFFC0000000000000000000" when X"32",
		X"FFFFFFFFFFFFE0000000000000000000" when X"33",
		X"FFFFFFFFFFFFF0000000000000000000" when X"34",
		X"FFFFFFFFFFFFF8000000000000000000" when X"35",
		X"FFFFFFFFFFFFFC000000000000000000" when X"36",
		X"FFFFFFFFFFFFFE000000000000000000" when X"37",
		X"FFFFFFFFFFFFFF000000000000000000" when X"38",
		X"FFFFFFFFFFFFFF800000000000000000" when X"39",
		X"FFFFFFFFFFFFFFC00000000000000000" when X"3A",
		X"FFFFFFFFFFFFFFE00000000000000000" when X"3B",
		X"FFFFFFFFFFFFFFF00000000000000000" when X"3C",
		X"FFFFFFFFFFFFFFF80000000000000000" when X"3D",
		X"FFFFFFFFFFFFFFFC0000000000000000" when X"3E",
		X"FFFFFFFFFFFFFFFE0000000000000000" when X"3F",
		X"FFFFFFFFFFFFFFFF0000000000000000" when X"40",
		X"FFFFFFFFFFFFFFFF8000000000000000" when X"41",
		X"FFFFFFFFFFFFFFFFC000000000000000" when X"42",
		X"FFFFFFFFFFFFFFFFE000000000000000" when X"43",
		X"FFFFFFFFFFFFFFFFF000000000000000" when X"44",
		X"FFFFFFFFFFFFFFFFF800000000000000" when X"45",
		X"FFFFFFFFFFFFFFFFFC00000000000000" when X"46",
		X"FFFFFFFFFFFFFFFFFE00000000000000" when X"47",
		X"FFFFFFFFFFFFFFFFFF00000000000000" when X"48",
		X"FFFFFFFFFFFFFFFFFF80000000000000" when X"49",
		X"FFFFFFFFFFFFFFFFFFC0000000000000" when X"4A",
		X"FFFFFFFFFFFFFFFFFFE0000000000000" when X"4B",
		X"FFFFFFFFFFFFFFFFFFF0000000000000" when X"4C",
		X"FFFFFFFFFFFFFFFFFFF8000000000000" when X"4D",
		X"FFFFFFFFFFFFFFFFFFFC000000000000" when X"4E",
		X"FFFFFFFFFFFFFFFFFFFE000000000000" when X"4F",
		X"FFFFFFFFFFFFFFFFFFFF000000000000" when X"50",
		X"FFFFFFFFFFFFFFFFFFFF800000000000" when X"51",
		X"FFFFFFFFFFFFFFFFFFFFC00000000000" when X"52",
		X"FFFFFFFFFFFFFFFFFFFFE00000000000" when X"53",
		X"FFFFFFFFFFFFFFFFFFFFF00000000000" when X"54",
		X"FFFFFFFFFFFFFFFFFFFFF80000000000" when X"55",
		X"FFFFFFFFFFFFFFFFFFFFFC0000000000" when X"56",
		X"FFFFFFFFFFFFFFFFFFFFFE0000000000" when X"57",
		X"FFFFFFFFFFFFFFFFFFFFFF0000000000" when X"58",
		X"FFFFFFFFFFFFFFFFFFFFFF8000000000" when X"59",
		X"FFFFFFFFFFFFFFFFFFFFFFC000000000" when X"5A",
		X"FFFFFFFFFFFFFFFFFFFFFFE000000000" when X"5B",
		X"FFFFFFFFFFFFFFFFFFFFFFF000000000" when X"5C",
		X"FFFFFFFFFFFFFFFFFFFFFFF800000000" when X"5D",
		X"FFFFFFFFFFFFFFFFFFFFFFFC00000000" when X"5E",
		X"FFFFFFFFFFFFFFFFFFFFFFFE00000000" when X"5F",
		X"FFFFFFFFFFFFFFFFFFFFFFFF00000000" when X"60",
		X"FFFFFFFFFFFFFFFFFFFFFFFF80000000" when X"61",
		X"FFFFFFFFFFFFFFFFFFFFFFFFC0000000" when X"62",
		X"FFFFFFFFFFFFFFFFFFFFFFFFE0000000" when X"63",
		X"FFFFFFFFFFFFFFFFFFFFFFFFF0000000" when X"64",
		X"FFFFFFFFFFFFFFFFFFFFFFFFF8000000" when X"65",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFC000000" when X"66",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFE000000" when X"67",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFF000000" when X"68",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFF800000" when X"69",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFFC00000" when X"6A",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFFE00000" when X"6B",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFFF00000" when X"6C",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFFF80000" when X"6D",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFFFC0000" when X"6E",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFFFE0000" when X"6F",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFFFF0000" when X"70",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFFFF8000" when X"71",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFC000" when X"72",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFE000" when X"73",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFF000" when X"74",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFF800" when X"75",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00" when X"76",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00" when X"77",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00" when X"78",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80" when X"79",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0" when X"7A",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0" when X"7B",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0" when X"7C",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8" when X"7D",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC" when X"7E",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE" when X"7F",
		X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF" when others;
end Behavioral;

